wait for 0.0000E+00 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='1';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 4.0000E-08 sec;
 MOSI<='0';
wait for 4.8000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 8.3860E-05 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.4000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 8.4300E-05 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='1';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 4.0000E-08 sec;
 MOSI<='0';
wait for 4.8000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 8.4280E-05 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 8.4280E-05 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 8.4300E-05 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 8.4300E-05 sec;
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.2000E-07 sec;
 SCK<='0';
wait for 4.8000E-07 sec;
 SCK<='1';
wait for 2.0000E-08 sec;
 MOSI<='0';
wait for 5.0000E-07 sec;
 SCK<='0';
wait for 5.0000E-07 sec;
 MOSI<='1';
 SCK<='1';
wait for 5.0000E-07 sec;
 SCK<='0';
